module online_adder_testing();

