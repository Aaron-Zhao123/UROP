library verilog;
use verilog.vl_types.all;
entity online_adder_testing is
    port(
        clk             : in     vl_logic
    );
end online_adder_testing;
