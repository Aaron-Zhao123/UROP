module four_bits_on_line_adder (x_plus,x_minus,y_plus,y_minus,clk,z_plus,z_minus);

	output[3:0] z_plus,z_minus;
	input clk;
	input [3:0] x_plus,x_minus,y_plus,y_minus;
	
	reg [5:0] z_plus_temp={}
	reg x_
	wire 
	
	